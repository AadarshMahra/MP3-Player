// top level 

