// top level 